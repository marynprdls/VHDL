library verilog;
use verilog.vl_types.all;
entity ejemplo1_vlg_vec_tst is
end ejemplo1_vlg_vec_tst;
